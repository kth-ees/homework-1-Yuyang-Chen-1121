module mul4(
    input logic [3:0] a,b,
    output logic [7:0] p
);
assign p = a*b;
endmodule
